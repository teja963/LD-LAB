module not_gate(b,a);
output b;
input a;
nand nand_1(b,a,a);
endmodule





