module not_gate_16(r,a);
output[15:0]r;
input[15:0]a;
not_gate not_gate_16[15:0](r,a);
endmodule


